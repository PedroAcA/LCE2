CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
30 0 30 100 9
65 72 715 758
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
59 Z:\home\paca\�rea de Trabalho\UnB\LCE2\CircuitMaker\BOM.DAT
0 7
65 72 715 758
144179219 0
0
6 Title:
5 Name:
0
0
0
14
10 Capacitor~
219 615 74 0 2 5
0 4 3
0
0 0 848 0
8 0.0708uF
-28 -18 28 -10
2 C4
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
8953 0 0
0
0
11 Signal Gen~
195 87 178 0 19 64
0 5 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 973279855
20
1 1000 0 0.0005 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
11 -500u/500uV
-39 -30 38 -22
2 V2
-7 -40 7 -32
0
0
39 %D %1 %2 DC 0 SIN(0 500u 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
4441 0 0
0
0
11 Signal Gen~
195 31 312 0 24 64
0 7 2 1 86 -10 10 0 0 0
0 0 0 0 0 0 0 1065353216 0 973279855
0 814313567 814313567 1056964608 1065353216
20
0 1 0 0.0005 0 1e-009 1e-009 0.5 1 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
7 0/500uV
-25 -30 24 -22
2 V1
-7 -40 7 -32
0
0
42 %D %1 %2 DC 0 PULSE(0 500u 0 1n 1n 500m 1)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3618 0 0
0
0
10 Capacitor~
219 153 297 0 2 5
0 6 2
0
0 0 848 0
5 100uF
-17 -18 18 -10
2 C3
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
6153 0 0
0
0
7 Ground~
168 238 372 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5394 0 0
0
0
7 Op Amp~
219 618 202 0 3 7
0 2 4 3
0
0 0 848 0
5 IDEAL
-18 -25 17 -17
2 U2
-7 -35 7 -27
0
0
17 %D %3 0 %1 %2 1E5
0
0
0
7

0 3 2 6 3 2 6 0
69 0 0 0 1 0 0 0
1 U
7734 0 0
0
0
7 Op Amp~
219 326 203 0 3 7
0 2 10 9
0
0 0 848 0
5 IDEAL
-18 -25 17 -17
2 U1
-7 -35 7 -27
0
0
17 %D %3 0 %1 %2 1E5
0
0
0
7

0 3 2 6 3 2 6 0
69 0 0 0 1 0 0 0
1 U
9914 0 0
0
0
10 Capacitor~
219 448 196 0 2 5
0 9 8
0
0 0 848 0
9 1.42857uF
-32 -18 31 -10
2 C2
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3747 0 0
0
0
10 Capacitor~
219 320 73 0 2 5
0 10 9
0
0 0 848 0
7 0.179uF
-25 -18 24 -10
2 C1
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3549 0 0
0
0
9 Resistor~
219 96 296 0 2 5
0 7 6
0
0 0 880 0
4 1.5k
-14 -14 14 -6
2 R5
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7931 0 0
0
0
9 Resistor~
219 616 143 0 2 5
0 4 3
0
0 0 880 0
6 561.9k
-21 -14 21 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9325 0 0
0
0
9 Resistor~
219 528 197 0 2 5
0 8 4
0
0 0 880 0
4 222k
-14 -14 14 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8903 0 0
0
0
9 Resistor~
219 323 144 0 2 5
0 10 9
0
0 0 880 0
4 220k
-14 -14 14 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3834 0 0
0
0
9 Resistor~
219 216 181 0 2 5
0 5 10
0
0 0 880 0
5 0.05k
-17 -14 18 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3363 0 0
0
0
20
2 0 3 0 0 8320 0 1 0 0 10 3
624 74
642 74
642 143
0 1 4 0 0 4224 0 0 1 11 0 3
588 143
588 74
606 74
2 0 2 0 0 12288 0 2 0 0 9 4
118 183
127 183
127 241
239 241
1 1 5 0 0 4224 0 2 14 0 0 4
118 173
190 173
190 181
198 181
0 0 2 0 0 0 0 0 0 6 20 2
170 314
238 314
2 2 2 0 0 0 0 3 4 0 0 5
62 317
62 330
170 330
170 297
162 297
2 1 6 0 0 12416 0 10 4 0 0 4
114 296
120 296
120 297
144 297
1 1 7 0 0 4224 0 3 10 0 0 4
62 307
75 307
75 296
78 296
1 0 2 0 0 0 0 7 0 0 20 3
308 209
239 209
239 300
2 3 3 0 0 0 0 11 6 0 0 4
634 143
644 143
644 202
636 202
0 1 4 0 0 0 0 0 11 12 0 3
585 197
585 143
598 143
2 2 4 0 0 0 0 12 6 0 0 4
546 197
592 197
592 196
600 196
2 1 8 0 0 4224 0 8 12 0 0 4
457 196
502 196
502 197
510 197
0 1 9 0 0 4224 0 0 8 15 0 2
352 196
439 196
0 3 9 0 0 0 0 0 7 16 0 4
349 144
352 144
352 203
344 203
2 2 9 0 0 0 0 9 13 0 0 4
329 73
349 73
349 144
341 144
0 1 10 0 0 8320 0 0 9 18 0 4
285 144
301 144
301 73
311 73
0 1 10 0 0 0 0 0 13 19 0 3
285 181
285 144
305 144
2 2 10 0 0 0 0 14 7 0 0 4
234 181
300 181
300 197
308 197
1 1 2 0 0 8320 0 6 5 0 0 4
600 208
600 300
238 300
238 366
0
0
8 0 0
0
0
0
0 0 0
0
0 0 0
100 0 0.001 4
0 5 0.01 0.01
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
655598 4356160 100 100 0 0
77 66 617 276
715 419 1365 767
523 66
77 66
617 135
617 276
0 0
3.30388 0.001 8057.14 0 3.999 3.999
12401 0
4 20 5000
1
644 178
0 3 0 0 2	0 10 0 0
590176 4356160 100 100 0 0
77 66 617 276
715 419 1365 767
602 66
77 66
617 275
617 276
0 0
5.53438e-315 5.26354e-315 5.2517e-315 0 5.53553e-315 5.53553e-315
12401 0
4 20 5000
1
564 169
0 5 0 0 2	0 10 0 0
983300 4356160 100 100 0 0
77 66 617 276
715 419 1365 767
617 66
77 66
617 263
617 276
0 0
0 0 0 0 0 0
12385 0
4 20 5000
1
644 153
0 6 0 0 2	0 10 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
